package apb_pkg;

import uvm_pkg::*;
`include "uvm_macros.svh"

`include "apb_transactions.svh"
`include "apb_scoreboard.svh"
`include "apb_sequences.svh"
`include "apb_monitor.svh"
`include "apb_driver.svh"
typedef uvm_sequencer#(apb_transaction) apb_sequencer;
`include "apb_agent.svh"
`include "apb_env.svh"
`include "apb_test.svh"

endpackage: apb_pkg
